//==============================================================================
// MAC Unit Module - Άσκηση 4
// Multiply and Accumulate Unit με 2 σειριακές ALUs
// Εκτελεί: result = (op1 * op2) + op3
//==============================================================================

module mac_unit (
    input  wire [31:0] op1,          // Πρώτη είσοδος (πολλαπλασιαστέος)
    input  wire [31:0] op2,          // Δεύτερη είσοδος (πολλαπλασιαστής/βάρος)
    input  wire [31:0] op3,          // Τρίτη είσοδος (πόλωση/bias)
    output wire [31:0] total_result, // Τελικό αποτέλεσμα MAC
    output wire        zero_mul,     // Ενεργό αν αποτέλεσμα πολ/σμού = 0
    output wire        zero_add,     // Ενεργό αν αποτέλεσμα πρόσθεσης = 0
    output wire        ovf_mul,      // Ενεργό αν υπερχείλιση στον πολ/σμό
    output wire        ovf_add       // Ενεργό αν υπερχείλιση στην πρόσθεση
);

    //--------------------------------------------------------------------------
    // Σταθερές για κωδικούς λειτουργίας ALU
    //--------------------------------------------------------------------------
    localparam [3:0] ALUOP_MULT = 4'b0110;  // Πολλαπλασιασμός
    localparam [3:0] ALUOP_ADD  = 4'b0100;  // Πρόσθεση

    //--------------------------------------------------------------------------
    // Ενδιάμεσα σήματα
    //--------------------------------------------------------------------------
    wire [31:0] mult_result;  // Αποτέλεσμα πολλαπλασιασμού

    //--------------------------------------------------------------------------
    // ALU 1: Πολλαπλασιασμός (op1 * op2)
    //--------------------------------------------------------------------------
    alu alu_mult (
        .op1    (op1),
        .op2    (op2),
        .alu_op (ALUOP_MULT),
        .zero   (zero_mul),
        .result (mult_result),
        .ovf    (ovf_mul)
    );

    //--------------------------------------------------------------------------
    // ALU 2: Πρόσθεση (mult_result + op3)
    //--------------------------------------------------------------------------
    alu alu_add (
        .op1    (mult_result),
        .op2    (op3),
        .alu_op (ALUOP_ADD),
        .zero   (zero_add),
        .result (total_result),
        .ovf    (ovf_add)
    );

endmodule

//==============================================================================
// Calculator Encoder Module - Άσκηση 2
// Structural Verilog - Παραγωγή alu_op από btnl, btnr, btnd
//
// Πίνακας Αλήθειας (από εκφώνηση):
// btnl btnr btnd | alu_op | Λειτουργία
// ----+----+----+---------+-----------
//  0    0    0  |  0000   | SRL
//  0    0    1  |  0101   | SLL
//  0    1    0  |  0100   | ADD
//  0    1    1  |  1100   | XOR
//  1    0    0  |  0010   | NOR
//  1    0    1  |  0111   | SUB
//  1    1    0  |  0110   | MULT
//  1    1    1  |  1111   | NAND
//
// Εξισώσεις από K-maps:
// alu_op[0] = btnd & (btnl | ~btnr)
// alu_op[1] = btnl
// alu_op[2] = btnr | btnd
// alu_op[3] = btnr & btnd
//==============================================================================

module calc_enc (
    input  wire btnl,           // Αριστερό πλήκτρο
    input  wire btnr,           // Δεξί πλήκτρο
    input  wire btnd,           // Κάτω πλήκτρο
    output wire [3:0] alu_op    // Κωδικός λειτουργίας ALU
);

    //--------------------------------------------------------------------------
    // Ενδιάμεσα σήματα
    //--------------------------------------------------------------------------
    wire btnr_n;                // NOT btnr
    wire or0_mid;               // btnl | (~btnr)

    //--------------------------------------------------------------------------
    // NOT πύλες - Σχ. 2
    //--------------------------------------------------------------------------
    not U_NOT_BTNR (btnr_n, btnr);

    //--------------------------------------------------------------------------
    // alu_op[0] = btnd & (btnl | ~btnr) - Σχ. 2
    // Πρώτα OR: btnl με ~btnr
    // Μετά AND: αποτέλεσμα με btnd
    //--------------------------------------------------------------------------
    or  U_OR0  (or0_mid, btnl, btnr_n);
    and U_AND0 (alu_op[0], btnd, or0_mid);

    //--------------------------------------------------------------------------
    // alu_op[1] = btnl - Σχ. 3
    // Απλή σύνδεση (buffer)
    //--------------------------------------------------------------------------
    buf U_BUF1 (alu_op[1], btnl);

    //--------------------------------------------------------------------------
    // alu_op[2] = btnr | btnd - Σχ. 4
    //--------------------------------------------------------------------------
    or U_OR2 (alu_op[2], btnr, btnd);

    //--------------------------------------------------------------------------
    // alu_op[3] = btnr & btnd - Σχ. 5
    //--------------------------------------------------------------------------
    and U_AND3 (alu_op[3], btnr, btnd);

endmodule

//==============================================================================
// ALU Module - Άσκηση 1
// 32-bit Arithmetic Logic Unit
//==============================================================================

module alu (
    input  wire [31:0] op1,      // Τελεστής 1 σε συμπλήρωμα ως προς 2
    input  wire [31:0] op2,      // Τελεστής 2 σε συμπλήρωμα ως προς 2
    input  wire [3:0]  alu_op,   // Κωδικός λειτουργίας
    output wire        zero,     // Ένδειξη μηδενικού αποτελέσματος
    output reg  [31:0] result,   // Αποτέλεσμα 32-bit
    output reg         ovf       // Ένδειξη υπερχείλισης
);

    //--------------------------------------------------------------------------
    // Ορισμός σταθερών για τους κωδικούς λειτουργίας της ALU
    //--------------------------------------------------------------------------
    parameter [3:0] ALUOP_AND   = 4'b1000;  // Λογική AND
    parameter [3:0] ALUOP_OR    = 4'b1001;  // Λογική OR
    parameter [3:0] ALUOP_NOR   = 4'b1010;  // Λογική NOR
    parameter [3:0] ALUOP_NAND  = 4'b1011;  // Λογική NAND
    parameter [3:0] ALUOP_XOR   = 4'b1100;  // Λογική XOR
    parameter [3:0] ALUOP_ADD   = 4'b0100;  // Προσημασμένη Πρόσθεση
    parameter [3:0] ALUOP_SUB   = 4'b0101;  // Προσημασμένη Αφαίρεση
    parameter [3:0] ALUOP_MULT  = 4'b0110;  // Προσημασμένος Πολλαπλασιασμός
    parameter [3:0] ALUOP_SRL   = 4'b0000;  // Λογική ολίσθηση δεξιά
    parameter [3:0] ALUOP_SLL   = 4'b0001;  // Λογική ολίσθηση αριστερά
    parameter [3:0] ALUOP_SRA   = 4'b0010;  // Αριθμητική ολίσθηση δεξιά
    parameter [3:0] ALUOP_SLA   = 4'b0011;  // Αριθμητική ολίσθηση αριστερά

    //--------------------------------------------------------------------------
    // Ενδιάμεσα σήματα για υπολογισμό υπερχείλισης
    //--------------------------------------------------------------------------
    wire [32:0] add_result;      // Αποτέλεσμα πρόσθεσης με επιπλέον bit
    wire [32:0] sub_result;      // Αποτέλεσμα αφαίρεσης με επιπλέον bit
    wire [63:0] mult_result;     // Πλήρες αποτέλεσμα πολλαπλασιασμού 64-bit
    
    // Επέκταση προσήμου για αριθμητικές πράξεις
    wire signed [31:0] op1_signed = op1;
    wire signed [31:0] op2_signed = op2;
    wire signed [63:0] mult_result_signed;
    
    // Υπολογισμός αποτελεσμάτων
    assign add_result = {op1[31], op1} + {op2[31], op2};
    assign sub_result = {op1[31], op1} - {op2[31], op2};
    assign mult_result_signed = op1_signed * op2_signed;
    assign mult_result = mult_result_signed;

    //--------------------------------------------------------------------------
    // Κύρια λογική ALU - Συνδυαστικό κύκλωμα
    //--------------------------------------------------------------------------
    always @(*) begin
        // Αρχικοποίηση εξόδων
        result = 32'b0;
        ovf = 1'b0;
        
        case (alu_op)
            //------------------------------------------------------------------
            // Λογικές πράξεις (χωρίς overflow)
            //------------------------------------------------------------------
            ALUOP_AND: begin
                result = op1 & op2;
                ovf = 1'b0;
            end
            
            ALUOP_OR: begin
                result = op1 | op2;
                ovf = 1'b0;
            end
            
            ALUOP_NOR: begin
                result = ~(op1 | op2);
                ovf = 1'b0;
            end
            
            ALUOP_NAND: begin
                result = ~(op1 & op2);
                ovf = 1'b0;
            end
            
            ALUOP_XOR: begin
                result = op1 ^ op2;
                ovf = 1'b0;
            end
            
            //------------------------------------------------------------------
            // Αριθμητικές πράξεις (με έλεγχο overflow)
            //------------------------------------------------------------------
            ALUOP_ADD: begin
                result = op1 + op2;
                // Overflow: αν τα πρόσημα των τελεστέων είναι ίδια και το πρόσημο
                // του αποτελέσματος διαφέρει
                ovf = (op1[31] == op2[31]) && (result[31] != op1[31]);
            end
            
            ALUOP_SUB: begin
                result = op1 - op2;
                // Overflow: αν τα πρόσημα διαφέρουν και το αποτέλεσμα έχει
                // το πρόσημο του op2
                ovf = (op1[31] != op2[31]) && (result[31] == op2[31]);
            end
            
            ALUOP_MULT: begin
                result = mult_result[31:0];
                // Overflow: αν τα υψηλότερα 33 bits δεν είναι όλα 0 ή όλα 1
                // (επέκταση προσήμου του bit 31)
                ovf = (mult_result[63:31] != {33{mult_result[31]}}) &&
                      (mult_result[63:31] != 33'b0);
            end
            
            //------------------------------------------------------------------
            // Πράξεις ολίσθησης (χωρίς overflow)
            //------------------------------------------------------------------
            ALUOP_SRL: begin  // Λογική ολίσθηση δεξιά
                result = op1 >> op2[4:0];  // Χρησιμοποιούμε μόνο τα 5 LSB του op2
                ovf = 1'b0;
            end
            
            ALUOP_SLL: begin  // Λογική ολίσθηση αριστερά
                result = op1 << op2[4:0];
                ovf = 1'b0;
            end
            
            ALUOP_SRA: begin  // Αριθμητική ολίσθηση δεξιά (διατηρεί πρόσημο)
                result = op1_signed >>> op2[4:0];
                ovf = 1'b0;
            end
            
            ALUOP_SLA: begin  // Αριθμητική ολίσθηση αριστερά
                result = op1_signed <<< op2[4:0];
                ovf = 1'b0;
            end
            
            default: begin
                result = 32'b0;
                ovf = 1'b0;
            end
        endcase
    end

    //--------------------------------------------------------------------------
    // Σήμα zero - ενεργό όταν το αποτέλεσμα είναι μηδέν
    //--------------------------------------------------------------------------
    assign zero = (result == 32'b0);

endmodule

//==============================================================================
// Calculator Testbench - Άσκηση 2
// Έλεγχος ορθής λειτουργίας αριθμομηχανής και ALU
//==============================================================================

`timescale 1ns / 1ps

module calc_tb;

    //--------------------------------------------------------------------------
    // Σήματα Testbench
    //--------------------------------------------------------------------------
    reg         clk;
    reg         btnc;
    reg         btnac;
    reg         btnl;
    reg         btnr;
    reg         btnd;
    reg  [15:0] sw;
    wire [15:0] led;
    
    // Μετρητής επιτυχών τεστ
    integer pass_count;
    integer test_count;

    //--------------------------------------------------------------------------
    // Instance του Calculator
    //--------------------------------------------------------------------------
    calc uut (
        .clk   (clk),
        .btnc  (btnc),
        .btnac (btnac),
        .btnl  (btnl),
        .btnr  (btnr),
        .btnd  (btnd),
        .sw    (sw),
        .led   (led)
    );

    //--------------------------------------------------------------------------
    // Δημιουργία σήματος ρολογιού - περίοδος 10ns
    //--------------------------------------------------------------------------
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    //--------------------------------------------------------------------------
    // Task για εκτέλεση πράξης στην αριθμομηχανή
    //--------------------------------------------------------------------------
    task execute_operation;
        input l, r, d;
        input [15:0] switch_val;
        input [15:0] expected;
        input [8*4-1:0] op_name; //Τα ονόματα των πράξεών έχουν έως 4 χαρακτήρες
        begin
            btnl = l;
            btnr = r;
            btnd = d;
            sw = switch_val;
            #1;  // Αναμονή για σταθεροποίηση σημάτων
            
            // Πάτημα κεντρικού πλήκτρου
            btnc = 1;
            @(posedge clk);
            #2;
            btnc = 0;
            #10;
            
            test_count = test_count + 1;
            
            // Έλεγχος αποτελέσματος
            if (led === expected) begin
                $display("PASS: %s - Expected: 0x%04h, Got: 0x%04h", 
                         op_name, expected, led);
                pass_count = pass_count + 1;
            end
            else begin
                $display("FAIL: %s - Expected: 0x%04h, Got: 0x%04h", 
                         op_name, expected, led);
            end
        end
    endtask

    //--------------------------------------------------------------------------
    // Task για reset
    //--------------------------------------------------------------------------
    task do_reset;
        begin
            btnac = 1;
            @(posedge clk);
            #2;
            btnac = 0;
            #10;
            
            test_count = test_count + 1;
            
            if (led === 16'h0000) begin
                $display("PASS: Reset - Expected: 0x0000, Got: 0x%04h", led);
                pass_count = pass_count + 1;
            end
            else begin
                $display("FAIL: Reset - Expected: 0x0000, Got: 0x%04h", led);
            end
        end
    endtask

    //--------------------------------------------------------------------------
    // Κύριο τεστ
    //--------------------------------------------------------------------------
    initial begin
        // Αρχικοποίηση
        $display("============================================================");
        $display("Calculator Testbench - Start");
        $display("============================================================");
        
        pass_count = 0;
        test_count = 0;
        btnc = 0;
        btnac = 0;
        btnl = 0;
        btnr = 0;
        btnd = 0;
        sw = 16'h0000;
        
        #20;
        
        //----------------------------------------------------------------------
        // Test 1: Reset (btnac)
        //----------------------------------------------------------------------
        $display("\n--- Test 1: Reset ---");
        do_reset();
        
        //----------------------------------------------------------------------
        // Test 2: ADD (btnl=0, btnr=1, btnd=0) -> alu_op = 0100
        // acc = 0x0 + 0x285a = 0x285a
        //----------------------------------------------------------------------
        $display("\n--- Test 2: ADD ---");
        execute_operation(0, 1, 0, 16'h285a, 16'h285a, "ADD");
        
        //----------------------------------------------------------------------
        // Test 3: XOR (btnl=1, btnr=1, btnd=1) -> alu_op = 1100
        // acc = 0x285a ^ 0x04c8 = 0x2c92
        //----------------------------------------------------------------------
        $display("\n--- Test 3: XOR ---");
        execute_operation(1, 1, 1, 16'h04c8, 16'h2c92, "XOR");
        
        //----------------------------------------------------------------------
        // Test 4: Logical Shift Right (btnl=0, btnr=0, btnd=0) -> alu_op = 0000
        // acc = 0x2c92 >> 5 = 0x0164
        //----------------------------------------------------------------------
        $display("\n--- Test 4: Logical Shift Right ---");
        execute_operation(0, 0, 0, 16'h0005, 16'h0164, "SRL");
        
        //----------------------------------------------------------------------
        // Test 5: NOR (btnl=1, btnr=0, btnd=1) -> alu_op = 1010
        // acc = ~(0x0164 | 0xa085) = 0x5e1a
        //----------------------------------------------------------------------
        $display("\n--- Test 5: NOR ---");
        execute_operation(1, 0, 1, 16'ha085, 16'h5e1a, "NOR");
        
        //----------------------------------------------------------------------
        // Test 6: MULT (btnl=1, btnr=0, btnd=0) -> alu_op = 0110
        // acc = 0x5e1a * 0x07fe = 0x2e74c (lower 16 bits = 0x13cc)
        // Σημείωση: 0x5e1a = 24090, 0x07fe = 2046
        // 24090 * 2046 = 49288140 = 0x2F013CC (16 LSB = 0x13CC)
        //----------------------------------------------------------------------
        $display("\n--- Test 6: MULT ---");
        execute_operation(1, 0, 0, 16'h07fe, 16'h13cc, "MULT");
        
        //----------------------------------------------------------------------
        // Test 7: Logical Shift Left (btnl=0, btnr=0, btnd=1) -> alu_op = 0001
        // acc = 0x13cc << 4 = 0x3cc0
        //----------------------------------------------------------------------
        $display("\n--- Test 7: Logical Shift Left ---");
        execute_operation(0, 0, 1, 16'h0004, 16'h3cc0, "SLL");
        
        //----------------------------------------------------------------------
        // Test 8: NAND (btnl=1, btnr=1, btnd=0) -> alu_op = 1011
        // acc = ~(0x3cc0 & 0xfa65) = ~(0x3840) = 0xc7bf
        //----------------------------------------------------------------------
        $display("\n--- Test 8: NAND ---");
        execute_operation(1, 1, 0, 16'hfa65, 16'hc7bf, "NAND");
        
        //----------------------------------------------------------------------
        // Test 9: SUB (btnl=0, btnr=1, btnd=1) -> alu_op = 0101
        // acc = 0xc7bf - 0xb2e4 = 0x14db
        // Σημείωση: 0xc7bf = -14401 (signed), 0xb2e4 = -19740 (signed)
        // -14401 - (-19740) = 5339 = 0x14DB
        //----------------------------------------------------------------------
        $display("\n--- Test 9: SUB ---");
        execute_operation(0, 1, 1, 16'hb2e4, 16'h14db, "SUB");
        
        //----------------------------------------------------------------------
        // Αποτελέσματα
        //----------------------------------------------------------------------
        $display("\n============================================================");
        $display("Calculator Testbench - Complete");
        $display("Results: %0d PASS / %0d Total Tests", pass_count, test_count);
        $display("============================================================");
        
        if (pass_count == test_count) begin
            $display("*** ALL TESTS PASSED ***");
        end
        else begin
            $display("*** SOME TESTS FAILED ***");
        end
        
        #100;
        $finish;
    end

    //--------------------------------------------------------------------------
    // Waveform dump για προσομοίωση
    //--------------------------------------------------------------------------
    initial begin
        $dumpfile("calc_tb.vcd");
        $dumpvars(0, calc_tb);
    end

endmodule

//==============================================================================
// Calculator Module - Άσκηση 2
// Αριθμομηχανή με accumulator 16-bit και ALU
//==============================================================================

module calc (
    input  wire        clk,     // Ρολόι
    input  wire        btnc,    // Κεντρικό πλήκτρο - εκτέλεση πράξης
    input  wire        btnac,   // Πλήκτρο εκκαθάρισης (all clear)
    input  wire        btnl,    // Αριστερό πλήκτρο
    input  wire        btnr,    // Δεξί πλήκτρο
    input  wire        btnd,    // Κάτω πλήκτρο
    input  wire [15:0] sw,      // Διακόπτες εισόδου δεδομένων
    output wire [15:0] led      // LED εξόδου του accumulator
);

    //--------------------------------------------------------------------------
    // Εσωτερικά σήματα
    //--------------------------------------------------------------------------
    reg  [15:0] accumulator;    // Καταχωρητής συσσωρευτή 16-bit
    wire [31:0] op1_extended;   // Επέκταση προσήμου του accumulator
    wire [31:0] op2_extended;   // Επέκταση προσήμου των switches
    wire [3:0]  alu_op;         // Κωδικός λειτουργίας ALU
    wire [31:0] alu_result;     // Αποτέλεσμα ALU
    wire        alu_zero;       // Σήμα zero της ALU
    wire        alu_ovf;        // Σήμα overflow της ALU

    //--------------------------------------------------------------------------
    // Επέκταση προσήμου (Sign Extension)
    // Επανάληψη του MSB για τα υψηλότερα 16 bits
    //--------------------------------------------------------------------------
    assign op1_extended = {{16{accumulator[15]}}, accumulator};
    assign op2_extended = {{16{sw[15]}}, sw};

    //--------------------------------------------------------------------------
    // Instance του ALU encoder (structural Verilog)
    //--------------------------------------------------------------------------
    calc_enc encoder_inst (
        .btnl   (btnl),
        .btnr   (btnr),
        .btnd   (btnd),
        .alu_op (alu_op)
    );

    //--------------------------------------------------------------------------
    // Instance της ALU
    //--------------------------------------------------------------------------
    alu alu_inst (
        .op1    (op1_extended),
        .op2    (op2_extended),
        .alu_op (alu_op),
        .zero   (alu_zero),
        .result (alu_result),
        .ovf    (alu_ovf)
    );

    //--------------------------------------------------------------------------
    // Καταχωρητής Accumulator
    // - Σύγχρονος μηδενισμός με btnac
    // - Ενημέρωση με btnc
    //--------------------------------------------------------------------------
    always @(posedge clk) begin
        if (btnac) begin
            // Σύγχρονος μηδενισμός
            accumulator <= 16'b0;
        end
        else if (btnc) begin
            // Ενημέρωση με τα 16 χαμηλότερα bits του αποτελέσματος
            accumulator <= alu_result[15:0];
        end
        // Αλλιώς διατήρηση της τρέχουσας τιμής
    end

    //--------------------------------------------------------------------------
    // Σύνδεση εξόδου LED με τον accumulator
    //--------------------------------------------------------------------------
    assign led = accumulator;

endmodule
